module decodetoBCD(
input in,
output[3:0]out1,out2);

reg  [7:0] out;

always @(*)
  case(in)
            6'b000000: out = 8'b00000000;//0
            
            6'b000001: out = 8'b00000001;
            6'b000010: out = 8'b00000010;
            6'b000011: out = 8'b00000011;
            6'b000100: out = 8'b00000100;
            6'b000101: out = 8'b00000101;
            6'b000110: out = 8'b00000110;
            6'b000111: out = 8'b00000111;
            6'b001000: out = 8'b00001000;
            6'b001001: out = 8'b00001001;
            
            6'b001010: out = 8'b00010000;//10
            
            6'b001011: out = 8'b00010001;
            6'b001100: out = 8'b00010010;
            6'b001101: out = 8'b00010011;
            6'b001110: out = 8'b00010100;
            6'b001111: out = 8'b00010101;
            6'b010000: out = 8'b00010110;
            6'b010001: out = 8'b00010111;
            6'b010010: out = 8'b00011000;
            6'b010011: out = 8'b00011001;
            
            6'b010100: out = 8'b00100000;//20
            
            6'b010101: out = 8'b00100001;
            6'b010110: out = 8'b00100010;
            6'b010111: out = 8'b00100011;
            6'b011000: out = 8'b00100100;
            6'b011001: out = 8'b00100101;
            6'b011010: out = 8'b00100110;
            6'b011011: out = 8'b00100111;
            6'b011100: out = 8'b00101000;
            6'b011101: out = 8'b00101001;
            
            6'b011110: out = 8'b00110000;//30
            
            6'b011111: out = 8'b00110001;
            6'b100000: out = 8'b00110010;
            6'b100001: out = 8'b00110011;
            6'b100010: out = 8'b00110100;
            6'b100011: out = 8'b00110101;
            6'b100100: out = 8'b00110110;
            6'b100101: out = 8'b00110111;
            6'b100110: out = 8'b00111000;
            6'b100111: out = 8'b00111001;
            
            6'b101000: out = 8'b01000000;//40
            
            6'b101001: out = 8'b01000001;
            6'b101010: out = 8'b01000010;
            6'b101011: out = 8'b01000011;
            6'b101100: out = 8'b01000100;
            6'b101101: out = 8'b01000101;
            6'b101110: out = 8'b01000110;
            6'b101111: out = 8'b01000111;
            6'b110000: out = 8'b01001000;
            6'b110001: out = 8'b01001001;
            
            6'b101000: out = 8'b01010000;//50
            
            6'b110010: out = 8'b01010001;
            6'b110011: out = 8'b01010010;
            6'b110100: out = 8'b01010011;
            6'b110101: out = 8'b01010100;
            6'b110110: out = 8'b01010101;
            6'b110111: out = 8'b01010110;
            6'b111000: out = 8'b01010111;
            6'b111001: out = 8'b01011000;
            6'b111010: out = 8'b01011001;
            
            6'b111100: out = 8'b01100000;//60
            
            default: out = 8'b00000000;
        endcase

assign {out2,out1} = out;

endmodule